----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:04:54 10/01/2020 
-- Design Name: 
-- Module Name:    ha_rtl - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ha_rtl is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
           carry : out  STD_LOGIC;
           sum : out  STD_LOGIC);
end ha_rtl;

architecture Behavioral of ha_rtl is

begin
	sum <= a xor b;
	carry <= a and b;

end Behavioral;

